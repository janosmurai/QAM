`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:53:40 03/23/2015 
// Design Name: 
// Module Name:    digit_BPS_filter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module digit_BPS_filter(
    input clock,
    input reset,
    input sgl_in,
    output sgl_out
    );


endmodule
