`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:26:42 03/23/2015 
// Design Name: 
// Module Name:    S2P 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module S2P(
    input clock,
    input reset,
    input adat_be_S,
    output  elojel_sin,
	 output  elojel_cos

    );


endmodule
